module axis_interconnect (
    ports
);
    
reg    [7:0] a;



    
end

endmodule